! This thermodynamic database was obtained by fitting the thermodynamic properties
! extracted from the following file: Thermodynamics.therm
! The thermodynamic properties are fitted in order to preserve not only the 
! continuity of each function at the intermediate temperature, but also the  continuity
! of the derivatives, from the 1st to the 3rd order
! The intermediate temperatures are the same for all the species.
! Last update: 12/22/2020

THERMO ALL
270.   1000.   3500. 
AR                      AR  1               G    200.00   3500.00 1000.00      1
 2.50020265e+00-5.42754143e-07 4.57710846e-10-1.53917542e-13 1.78608595e-17    2
-7.45429770e+02 4.37863370e+00 2.49980451e+00 1.04980652e-06-1.93113014e-09    3
 1.43864312e-12-3.80279305e-16-7.45350142e+02 4.38055449e+00                   4
N2                      N   2               G    200.00   3500.00 1000.00      1
 2.86705237e+00 1.54614237e-03-5.84320220e-07 1.02525351e-10-6.87117090e-15    2
-8.88091985e+02 6.35154244e+00 3.75165514e+00-1.99226869e-03 4.72329636e-06    3
-3.43588570e-09 8.77731593e-13-1.06501254e+03 2.08384546e+00                   4
HE                      HE  1               G    200.00   3500.00 1000.00      1
 2.50028359e+00-7.18471398e-07 5.99685721e-10-2.00458035e-13 2.31417158e-17    2
-7.45453089e+02 9.27233751e-01 2.49971505e+00 1.55569518e-06-2.81156415e-09    3
 2.07370855e-12-5.45399930e-16-7.45339381e+02 9.29976636e-01                   4
H2                      H   2               G    200.00   3500.00 1000.00      1
 3.97161381e+00-1.44148688e-03 1.56248342e-06-5.19085786e-10 5.86218466e-14    2
-1.16573011e+03-6.62288576e+00 3.03115666e+00 2.32034174e-03-4.08025952e-06    3
 3.24274284e-09-8.81835310e-13-9.77638676e+02-2.08572362e+00                   4
H                       H   1               G    200.00   3500.00 1000.00      1
 2.50042553e+00-1.02575684e-06 8.34881465e-10-2.74914263e-13 3.14676920e-17    2
 2.54736098e+04-4.48949941e-01 2.49959101e+00 2.31230761e-06-4.17221522e-09    3
 3.06315020e-12-8.03048423e-16 2.54737767e+04-4.44923883e-01                   4
O2                      O   2               G    200.00   3500.00 1000.00      1
 2.65938544e+00 2.84309875e-03-1.78721131e-06 5.35030074e-10-5.83386805e-14    2
-8.76533747e+02 8.81275457e+00 3.43324602e+00-2.52343589e-04 2.85595221e-06    3
-2.56041227e-09 7.15521905e-13-1.03130586e+03 5.07932458e+00                   4
O                       O   1               G    200.00   3500.00 1000.00      1
 2.50518318e+00 7.18274073e-05-8.72697956e-08 3.28327158e-11-3.72698409e-15    2
 2.92429404e+04 5.12195346e+00 3.00862935e+00-1.94195728e-03 2.93340724e-06    3
-1.98095197e-09 4.99719188e-13 2.91422512e+04 2.69311670e+00                   4
H2O                     H   2O   1          G    200.00   3500.00 1000.00      1
 3.33911324e+00 1.65341899e-03 1.25490864e-07-1.70489006e-10 2.41757907e-14    2
-3.01285262e+04 3.26058181e+00 4.16994328e+00-1.66990116e-03 5.11047110e-06    3
-3.49380916e-09 8.55005830e-13-3.02946923e+04-7.47692860e-01                   4
OH                      H   1O   1          G    200.00   3500.00 1000.00      1
 3.54142511e+00-4.02539504e-04 8.28983436e-07-3.06007231e-10 3.59487658e-14    2
 3.47772231e+03 2.04510885e+00 3.97872055e+00-2.15172124e-03 3.45275604e-06    3
-2.05518897e-09 4.73244200e-13 3.39026323e+03-6.45888421e-02                   4
H2O2                    H   2O   2          G    200.00   3500.00 1000.00      1
 3.51570577e+00 6.39707142e-03-2.99616894e-06 7.29517164e-10-7.03368251e-14    2
-1.76035639e+04 6.37746731e+00 3.37185986e+00 6.97245505e-03-3.85924438e-06    3
 1.30490079e-09-2.14182732e-13-1.75747947e+04 7.07144066e+00                   4
HO2                     H   1O   2          G    200.00   3500.00 1000.00      1
 3.03708588e+00 4.39299607e-03-2.14979388e-06 5.79665495e-10-6.20606503e-14    2
 4.02463864e+02 9.05743987e+00 3.34368647e+00 3.16659373e-03-3.10190367e-07    3
-6.46736847e-10 2.44539935e-13 3.41143747e+02 7.57826927e+00                   4
NO                      N   1O   1          G    200.00   3500.00 1000.00      1
 2.59354221e+00 2.64415882e-03-1.52114885e-06 4.10403638e-10-4.18254553e-14    2
 1.01483561e+04 9.96631515e+00 4.01174047e+00-3.02863423e-03 6.98804072e-06    3
-5.26238941e-09 1.37637281e-12 9.86471645e+03 3.12432834e+00                   4
N2O                     N   2O   1          G    200.00   3500.00 1000.00      1
 3.73479467e+00 4.92112867e-03-2.64141082e-06 6.75979379e-10-6.61701157e-14    2
 8.45788435e+03 3.70529413e+00 2.32814393e+00 1.05477316e-02-1.10813152e-05    3
 6.30258232e-09-1.47282085e-12 8.73921450e+03 1.04915708e+01                   4
NO2                     N   1O   2          G    200.00   3500.00 1000.00      1
 2.81928760e+00 6.66768363e-03-4.20601408e-06 1.21236128e-09-1.27472160e-13    2
 3.01997287e+03 1.10216156e+01 3.02085906e+00 5.86139777e-03-2.99658531e-06    3
 4.06075432e-10 7.40993029e-14 2.97965858e+03 1.00491498e+01                   4
HNO                     H   1N   1O   1     G    200.00   3500.00 1000.00      1
 2.58538362e+00 4.39768557e-03-1.51527792e-06 3.27344483e-10-3.48008773e-14    2
 1.19447198e+04 1.07066015e+01 3.95390792e+00-1.07641160e-03 6.69586784e-06    3
-5.14675269e-09 1.33372342e-12 1.16710149e+04 4.10426287e+00                   4
HNO2                    H   1N   1O   2     G    200.00   3500.00 1000.00      1
 1.67672720e+00 1.13742369e-02-6.65140747e-06 1.80801424e-09-1.85461497e-13    2
-6.22986791e+03 1.60907952e+01 2.50761895e+00 8.05066991e-03-1.66605697e-06    3
-1.51555276e-09 6.45430253e-13-6.39604626e+03 1.20822228e+01                   4
HONO                    H   1N   1O   2     G    200.00   3500.00 1000.00      1
 4.27918633e+00 6.88970202e-03-3.70392984e-06 9.54587536e-10-9.47191408e-14    2
-1.10731255e+04 4.10913869e+00 2.48864620e+00 1.40518625e-02-1.44471706e-05    3
 8.11674804e-09-1.88525927e-12-1.07150175e+04 1.27474598e+01                   4
HONO2                   H   1N   1O   3     G    200.00   3500.00 1000.00      1
 4.53382238e+00 1.19894623e-02-7.32618265e-06 2.02955283e-09-2.09762347e-13    2
-1.81055423e+04 2.64544358e+00 6.03055389e-01 2.77125303e-02-3.09107846e-05    3
 1.77526208e-08-4.14052934e-12-1.73193889e+04 2.16091221e+01                   4
N2H2                    N   2H   2          G    300.00   3500.00 1000.00      1
 1.97737018e+00 8.91844494e-03-4.40431229e-06 1.05190934e-09-9.80620109e-14    2
 2.42198218e+04 1.25741464e+01 2.48823124e+00 6.87500070e-03-1.33914593e-06    3
-9.91534900e-10 4.12799049e-13 2.41176496e+04 1.01095371e+01                   4
H2NN                    N   2H   2          G    200.00   3500.00 1000.00      1
 9.69068217e-01 1.07127806e-02-5.61487273e-06 1.41593821e-09-1.38510047e-13    2
 3.55686201e+04 1.79803472e+01 3.60942403e+00 1.51357329e-04 1.02272621e-05    3
-9.14548503e-09 2.50184576e-12 3.50405489e+04 5.24215669e+00                   4
NH2OH                   N   1H   3O   1     G    200.00   3500.00 1000.00      1
 3.62592572e+00 8.71790060e-03-3.25468337e-06 5.74069573e-10-4.06039679e-14    2
-6.77351878e+03 5.16631665e+00 2.29706787e+00 1.40333320e-02-1.12278305e-05    3
 5.88950100e-09-1.36946183e-12-6.50774721e+03 1.15772877e+01                   4
HNOH                    H   2N   1O   1     G    200.00   3500.00 1000.00      1
 2.58923565e+00 7.95626702e-03-3.97699932e-06 9.87009095e-10-9.64164196e-14    2
 1.10468780e+04 1.11269069e+01 2.67978764e+00 7.59405907e-03-3.43368741e-06    3
 6.24801150e-10-5.86443340e-15 1.10287676e+04 1.06900459e+01                   4
NH3                     H   3N   1          G    200.00   3500.00 1000.00      1
 2.17000818e+00 6.76363558e-03-2.64200998e-06 5.26178719e-10-4.21542607e-14    2
-6.35633825e+03 9.03526090e+00 3.58776922e+00 1.09259142e-03 5.86455626e-06    3
-5.14486544e-09 1.37560678e-12-6.63989046e+03 2.19538342e+00                   4
N2H4                    N   2H   4          G    200.00   3500.00 1000.00      1
 2.51016628e+00 1.40719894e-02-7.01651081e-06 1.72966000e-09-1.67845607e-13    2
 1.01045064e+04 1.03911368e+01 1.66158577e+00 1.74663115e-02-1.21079939e-05    3
 5.12398203e-09-1.01642612e-12 1.02742225e+04 1.44850472e+01                   4
N                       N   1               G    200.00   3500.00 1000.00      1
 2.49388718e+00 1.03463894e-05 1.86373408e-09-6.88831040e-12 2.02531947e-15    2
 5.61062734e+04 4.22664618e+00 2.50529382e+00-3.52801814e-05 7.03035902e-08    3
-5.25148812e-11 1.34319622e-14 5.61039921e+04 4.17161573e+00                   4
NO3                     N   1O   3          G    200.00   3500.00 1000.00      1
 4.63338302e+00 8.75778392e-03-5.64510346e-06 1.61870163e-09-1.71019250e-13    2
 7.10564604e+03 1.22164434e+00 2.83089005e-01 2.61589600e-02-3.17468676e-05    3
 1.90198777e-08-4.52131327e-12 7.97570484e+03 2.22092983e+01                   4
NH                      N   1H   1          G    200.00   3500.00 1000.00      1
 3.35042867e+00 7.69077379e-05 5.26498857e-07-2.20844533e-10 2.78392313e-14    2
 4.21570028e+04 2.69491259e+00 3.70661261e+00-1.34782800e-03 2.66360247e-06    3
-1.64558027e-09 3.84023166e-13 4.20857660e+04 9.76530994e-01                   4
NNH                     N   2H   1          G    200.00   3500.00 1000.00      1
 2.37841845e+00 5.49090820e-03-2.85625537e-06 7.13106252e-10-6.91355603e-14    2
 2.91296358e+04 1.20624183e+01 3.89754146e+00-5.85583840e-04 6.25848270e-06    3
-5.36338579e-09 1.44998745e-12 2.88258112e+04 4.73352793e+00                   4
NH2                     N   1H   2          G    200.00   3500.00 1000.00      1
 3.07029783e+00 2.43321667e-03-2.97441803e-07-9.59510694e-11 2.14387823e-14    2
 2.14120013e+04 5.33199326e+00 4.22292679e+00-2.17729917e-03 6.61833196e-06    3
-4.70646691e-09 1.17406774e-12 2.11814755e+04-2.28775188e-01                   4
H2NO                    N   1H   2O   1     G    200.00   3500.00 1000.00      1
 2.60469506e+00 7.67251442e-03-3.65359694e-06 8.66020061e-10-8.16618809e-14    2
 6.90925077e+03 1.05131689e+01 3.32193214e+00 4.80356610e-03 6.49825548e-07    3
-2.00292826e-09 6.35575200e-13 6.76580336e+03 7.05291457e+00                   4
N2H3                    N   2H   3          G    200.00   3500.00 1000.00      1
 2.44355092e+00 1.08055013e-02-5.10970944e-06 1.20836975e-09-1.13960343e-13    2
 2.58683149e+04 1.15160769e+01 2.13725406e+00 1.20306887e-02-6.94749058e-06    3
 2.43355717e-09-4.20257198e-13 2.59295743e+04 1.29937821e+01                   4
END
